module part9()

endmodule
