module part3(input [7:0]SW,
				 input [2:1]KEY,
				 input CLOCK_50,
				 output [6:0]HEX0,
				 output [6:0]HEX1,
				 output [6:0]HEX2);
	wire [7:0]count;
	wire [3:0]bcd0,bcd1,bcd2;
	wire [11:0]counter;
	wire enable;
				 
	Clock_divider toSec(CLOCK_50,32'd50000000,CLOCK_sec);
	Clock_divider toMSec(CLOCK_50,32'd50000,CLOCK_msec);
	secCount count1(SW[7:0],CLOCK_sec,KEY[1],enable,count);
	msecCount count2(CLOCK_msec,KEY[1],enable,KEY[2],counter[11:0]);
	
	BintoBCD converter(counter,bcd0[3:0],bcd1[3:0],bcd2[3:0]);
	BCDto7 hex0(bcd0,HEX0);
	BCDto7 hex1(bcd1,HEX1);
	BCDto7 hex2(bcd2,HEX2);
				 
endmodule 

module BCDto7(input [3:0]sw,
				 output [6:0]hex);
				 
	assign hex[0] =  ~(sw[3] | sw[1] | (sw[2] ~^ sw[0]));
	assign hex[1] =  ~(~sw[2] | (sw[0] ~^ sw[1]));
	assign hex[2] =  ~(sw[2] | ~sw[1] | sw[0]);
	assign hex[3] =  ~(~sw[2]&~sw[0] | sw[1]&~sw[0] | sw[2]&~sw[1]&sw[0] | ~sw[2]&sw[1] | sw[3]);
	assign hex[4] =  ~(~sw[2]&~sw[0] | sw[1]&~sw[0]);
	assign hex[5] =  ~(sw[3] | ~sw[1]&~sw[0] | sw[2]&~sw[1] | sw[2]&~sw[0]);
	assign hex[6] =  ~(sw[3] | sw[1]&~sw[0] | sw[2]^sw[1]);
	
endmodule

module BintoBCD(input [11:0]bin,
					 output [3:0]bcd0,bcd1,bcd2);
			
	assign bcd0 = bin%7'd10;
	assign bcd1 = (bin/7'd10)%10;
	assign bcd2 = bin/100;
endmodule

module Clock_divider(input clock_in,
							input [31:0]DIVISOR,
							output reg clock_out);

	reg[31:0] counter=32'd0;
	
	always @(posedge clock_in)
	begin
		counter <= counter + 32'd1;
		if(counter>=(DIVISOR-1))
			counter <= 32'd0;
	end

	//assign clock_out = (counter<DIVISOR/2)?1'b0:1'b1;
	always@(posedge clock_in)
	begin
		if (counter<DIVISOR/2)
			clock_out = 1'b0;
		else 
			clock_out = 1'b1;
	end
endmodule

module secCount(input [7:0]load,
					 input ClkS,
					 input reset,
					 output rollOver,
					 output reg [7:0]countSec);

	//reg [7:0]countSec;	
					
	always@(posedge ClkS or negedge reset)
	begin
		if (reset == 0)
		begin
			countSec <= load;
		end
		
		else
		begin
			if (countSec == 0)
				countSec <= countSec;
			else
				countSec <= countSec - 1'b1;
		end
	end
	
	assign rollOver = (countSec == 0)? 1'b1:1'b0;
					 
endmodule

module msecCount(input ClkMS,
					  input reset,
					  input enable,
					  input stop,
					  output reg [11:0]countmSec);

	reg increment;
	
	always@(posedge ClkMS or negedge stop or negedge reset)
		begin
			if (reset == 0)
			begin
					countmSec <= 1'b0;
					increment <= 1;
			end
			else if(!stop)
				increment <= 0 | ~enable;
			else if (enable == 1)
				countmSec <= countmSec + increment;
		end
endmodule

module tb();
	reg CLOCK_50;
	reg [7:0]sw;
	reg reset,reaction;
	wire [6:0]hex0,hex1,hex2;
	wire [7:0]count;
	wire clkms, clks;
	
	
	
	part3 test(sw[7:0],{reaction,reset},CLOCK_50,hex0,hex1,hex2,count);
	
	
	assign clkms = test.CLOCK_msec;
	assign clks = test.CLOCK_sec;
	
	initial begin
		#0 	CLOCK_50 = 1'b0; 	sw = 8'd20;	reset = 1;	reaction = 1;
		#100 	CLOCK_50 = 1'b1;	reset = 0;
		#100 	CLOCK_50 = 1'b0;	reset = 0;
		#100 	CLOCK_50 = 1'b1;	reset = 0;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;	reset = 1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;	
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;	reaction = 0;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;	reaction = 1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		#100 	CLOCK_50 = 1'b0;
		#100 	CLOCK_50 = 1'b1;
		
	end
endmodule