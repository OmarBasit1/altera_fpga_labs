module part4()

endmodule 