module part3()
	
endmodule