module part7();

endmodule

// miss