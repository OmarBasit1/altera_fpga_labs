module part2()

endmodule

//same as in part 1